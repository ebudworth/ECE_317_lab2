i   �������?���ư>                �� B`��"۹?�������?���ư>      �?                                    @2                 V1      V1 �    �   �      )\���(�?      @	           6                 VP1     I01 ��� �  �   	           6                 VP2  W I02 W �   �      ���מYB?2                  L1 �����L1 �      �              -C��6?2                 C1  i r C1  o u @  �                     9@2                 R1     R1     `  �                      �      �   �   �   �                              �      �   �   �   �                              �   	   (  �   @  �                              �   
   @  �   `  �                              �      `  �   �  �                              �      `    �                               �      @    `                               �      �     @                               �      �     �                                �                 GND1 ��� ���    �        